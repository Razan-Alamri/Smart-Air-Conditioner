<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-49.2175,45.6776,58.6775,-7.91556</PageViewport>
<gate>
<ID>1</ID>
<type>AA_TOGGLE</type>
<position>-48,35</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>-48,39</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>DE_TO</type>
<position>-43.5,35</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Timer</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>-15,18</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-48,31</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>-40.5,31</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>-42,28.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>-28.5,15</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Timer</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_AND2</type>
<position>-4.5,15</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-48,43</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>8,17</position>
<gparam>LABEL_TEXT D</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-43.5,43</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Temperature Sensor</lparam></gate>
<gate>
<ID>33</ID>
<type>AE_DFF_LOW</type>
<position>12,13</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUTINV_0</ID>35 </output>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clear</ID>49 </input>
<input>
<ID>clock</ID>36 </input>
<input>
<ID>set</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>34</ID>
<type>DE_TO</type>
<position>-43.5,39</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Motion Sensor</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>9,29</position>
<gparam>LABEL_TEXT High Temperature</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>10,1</position>
<gparam>LABEL_TEXT Low Temperature</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>-43.5,31</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>40</ID>
<type>DA_FROM</type>
<position>-28,21</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Motion Sensor</lparam></gate>
<gate>
<ID>42</ID>
<type>DA_FROM</type>
<position>-20,9</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>37,4</position>
<gparam>LABEL_TEXT Razan Alamri</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>36.5,1</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>36,-2</position>
<gparam>LABEL_TEXT CAR</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>-6,26</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Temperature Sensor</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>26,17</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>26,10</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>BB_CLOCK</type>
<position>-3,8.5</position>
<output>
<ID>CLK</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>34.5,10.5</position>
<gparam>LABEL_TEXT A/C OFF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>33.5,17.5</position>
<gparam>LABEL_TEXT A/C ON</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-46,35,-45.5,35</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<connection>
<GID>3</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,21,-22,21</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>-22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-22,19,-22,21</points>
<intersection>19 4</intersection>
<intersection>21 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-22,19,-18,19</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>-22 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,15,-22,17</points>
<intersection>15 2</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-22,17,-18,17</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,15,-22,15</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-22 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1.5,15,9,15</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-46,31,-45.5,31</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,9,-12,14</points>
<intersection>9 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,14,-7.5,14</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-18,9,-12,9</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,16,-12,18</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12,16,-7.5,16</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-12 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,43,-45.5,43</points>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-46,39,-45.5,39</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,15,20,17</points>
<intersection>15 2</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,17,25,17</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,15,20,15</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,10,20,12</points>
<intersection>10 1</intersection>
<intersection>12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,10,25,10</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,12,20,12</points>
<connection>
<GID>33</GID>
<name>OUTINV_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4,8.5,4,12</points>
<intersection>8.5 2</intersection>
<intersection>12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,12,9,12</points>
<connection>
<GID>33</GID>
<name>clock</name></connection>
<intersection>4 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,8.5,4,8.5</points>
<connection>
<GID>56</GID>
<name>CLK</name></connection>
<intersection>4 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,3,6,26</points>
<intersection>3 3</intersection>
<intersection>26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,26,12,26</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>6 0</intersection>
<intersection>12 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>6,3,12,3</points>
<intersection>6 0</intersection>
<intersection>12 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>12,17,12,26</points>
<connection>
<GID>33</GID>
<name>set</name></connection>
<intersection>26 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>12,3,12,9</points>
<connection>
<GID>33</GID>
<name>clear</name></connection>
<intersection>3 3</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>31.6407,-2.39329,175.501,-73.851</PageViewport>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>46,-42.5</position>
<gparam>LABEL_TEXT </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>BA_NAND2</type>
<position>102.5,-19.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>BA_NAND2</type>
<position>102.5,-44.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>BA_NAND2</type>
<position>127.5,-26.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>127.5,-37.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>145,-37.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>145,-26.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>HE_JUNC_4</type>
<position>134.5,-37.5</position>
<input>
<ID>N_in0</ID>39 </input>
<input>
<ID>N_in1</ID>40 </input>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>HE_JUNC_4</type>
<position>134.5,-26.5</position>
<input>
<ID>N_in0</ID>42 </input>
<input>
<ID>N_in1</ID>41 </input>
<input>
<ID>N_in2</ID>44 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>95.5,-18.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Temperaturr>22</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>94.5,-45.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Temperaturr22</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>150.5,-37</position>
<gparam>LABEL_TEXT OFF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>150,-26</position>
<gparam>LABEL_TEXT ON</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AE_OR2</type>
<position>75.5,-36</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>65.5,-32</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Motion Sensor</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>65.5,-40</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>84</ID>
<type>DA_FROM</type>
<position>75,-42</position>
<input>
<ID>IN_0</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Control</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>88,-37</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115.5,-25.5,115.5,-19.5</points>
<intersection>-25.5 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115.5,-25.5,124.5,-25.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>115.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>105.5,-19.5,115.5,-19.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>115.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114.5,-44.5,114.5,-38.5</points>
<intersection>-44.5 1</intersection>
<intersection>-38.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105.5,-44.5,114.5,-44.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>114.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>114.5,-38.5,124.5,-38.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>114.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130.5,-37.5,133.5,-37.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-37.5,144,-37.5</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<connection>
<GID>73</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-26.5,144,-26.5</points>
<connection>
<GID>76</GID>
<name>N_in1</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130.5,-26.5,133.5,-26.5</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-32.5,121.5,-27.5</points>
<intersection>-32.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-27.5,124.5,-27.5</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-32.5,134.5,-32.5</points>
<intersection>121.5 0</intersection>
<intersection>134.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>134.5,-36.5,134.5,-32.5</points>
<connection>
<GID>75</GID>
<name>N_in3</name></connection>
<intersection>-32.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-31.5,134.5,-27.5</points>
<connection>
<GID>76</GID>
<name>N_in2</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-31.5,134.5,-31.5</points>
<intersection>122.5 2</intersection>
<intersection>134.5 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>122.5,-36.5,122.5,-31.5</points>
<intersection>-36.5 3</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>122.5,-36.5,124.5,-36.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>122.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-43.5,96.5,-20.5</points>
<intersection>-43.5 1</intersection>
<intersection>-37 4</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-43.5,99.5,-43.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>96.5,-20.5,99.5,-20.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>91,-37,96.5,-37</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,-18.5,99.5,-18.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>96.5,-45.5,99.5,-45.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-35,70.5,-32</points>
<intersection>-35 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-32,70.5,-32</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-35,72.5,-35</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-40,70.5,-37</points>
<intersection>-40 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-40,70.5,-40</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-37,72.5,-37</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78.5,-36,85,-36</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-42,80.5,-38</points>
<intersection>-42 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-38,85,-38</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-42,80.5,-42</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 2>
<page 3>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 3>
<page 4>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 4>
<page 5>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 5>
<page 6>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 6>
<page 7>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 7>
<page 8>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 8>
<page 9>
<PageViewport>-24.3048,25.3499,231.447,-101.686</PageViewport></page 9></circuit>